/run/media/user1/c2s/sriram/SCLPDK/scl_pdk/iolib/cio150/cds/lef/tsl18cio150_4lm.lef