/run/media/user1/c2s/sriram/SCLPDK/scl_pdk/stdlib/fs120/tech_data/lef/tsl180l4.lef